module add1(input [47:0]a, output [47:0]b);
assign b=a + 1'b1;
endmodule
